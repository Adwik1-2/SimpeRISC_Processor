module lsl(
    input  [31:0] d,         // Input data
    input  [4:0]  sel,       // Shift amount (0–31)
    output [31:0] y          // Output after logical left shift
);
    wire [31:0] stage1, stage2, stage3, stage4, stage5;

    // Shift by 1 if sel[0] is set
    assign stage1[0]  = sel[0] ? d[1]  : d[0];
    assign stage1[1]  = sel[0] ? d[2]  : d[1];
    assign stage1[2]  = sel[0] ? d[3]  : d[2];
    assign stage1[3]  = sel[0] ? d[4]  : d[3];
    assign stage1[4]  = sel[0] ? d[5]  : d[4];
    assign stage1[5]  = sel[0] ? d[6]  : d[5];
    assign stage1[6]  = sel[0] ? d[7]  : d[6];
    assign stage1[7]  = sel[0] ? d[8]  : d[7];
    assign stage1[8]  = sel[0] ? d[9]  : d[8];
    assign stage1[9]  = sel[0] ? d[10] : d[9];
    assign stage1[10] = sel[0] ? d[11] : d[10];
    assign stage1[11] = sel[0] ? d[12] : d[11];
    assign stage1[12] = sel[0] ? d[13] : d[12];
    assign stage1[13] = sel[0] ? d[14] : d[13];
    assign stage1[14] = sel[0] ? d[15] : d[14];
    assign stage1[15] = sel[0] ? d[16] : d[15];
    assign stage1[16] = sel[0] ? d[17] : d[16];
    assign stage1[17] = sel[0] ? d[18] : d[17];
    assign stage1[18] = sel[0] ? d[19] : d[18];
    assign stage1[19] = sel[0] ? d[20] : d[19];
    assign stage1[20] = sel[0] ? d[21] : d[20];
    assign stage1[21] = sel[0] ? d[22] : d[21];
    assign stage1[22] = sel[0] ? d[23] : d[22];
    assign stage1[23] = sel[0] ? d[24] : d[23];
    assign stage1[24] = sel[0] ? d[25] : d[24];
    assign stage1[25] = sel[0] ? d[26] : d[25];
    assign stage1[26] = sel[0] ? d[27] : d[26];
    assign stage1[27] = sel[0] ? d[28] : d[27];
    assign stage1[28] = sel[0] ? d[29] : d[28];
    assign stage1[29] = sel[0] ? d[30] : d[29];
    assign stage1[30] = sel[0] ? d[31] : d[30];
    assign stage1[31] = sel[0] ? 1'b0  : d[31];   // LSB shifted in as 0

    // Shift by 2 if sel[1] is set
    assign stage2[0]  = sel[1] ? stage1[2]  : stage1[0];
    assign stage2[1]  = sel[1] ? stage1[3]  : stage1[1];
    assign stage2[2]  = sel[1] ? stage1[4]  : stage1[2];
    assign stage2[3]  = sel[1] ? stage1[5]  : stage1[3];
    assign stage2[4]  = sel[1] ? stage1[6]  : stage1[4];
    assign stage2[5]  = sel[1] ? stage1[7]  : stage1[5];
    assign stage2[6]  = sel[1] ? stage1[8]  : stage1[6];
    assign stage2[7]  = sel[1] ? stage1[9]  : stage1[7];
    assign stage2[8]  = sel[1] ? stage1[10] : stage1[8];
    assign stage2[9]  = sel[1] ? stage1[11] : stage1[9];
    assign stage2[10] = sel[1] ? stage1[12] : stage1[10];
    assign stage2[11] = sel[1] ? stage1[13] : stage1[11];
    assign stage2[12] = sel[1] ? stage1[14] : stage1[12];
    assign stage2[13] = sel[1] ? stage1[15] : stage1[13];
    assign stage2[14] = sel[1] ? stage1[16] : stage1[14];
    assign stage2[15] = sel[1] ? stage1[17] : stage1[15];
    assign stage2[16] = sel[1] ? stage1[18] : stage1[16];
    assign stage2[17] = sel[1] ? stage1[19] : stage1[17];
    assign stage2[18] = sel[1] ? stage1[20] : stage1[18];
    assign stage2[19] = sel[1] ? stage1[21] : stage1[19];
    assign stage2[20] = sel[1] ? stage1[22] : stage1[20];
    assign stage2[21] = sel[1] ? stage1[23] : stage1[21];
    assign stage2[22] = sel[1] ? stage1[24] : stage1[22];
    assign stage2[23] = sel[1] ? stage1[25] : stage1[23];
    assign stage2[24] = sel[1] ? stage1[26] : stage1[24];
    assign stage2[25] = sel[1] ? stage1[27] : stage1[25];
    assign stage2[26] = sel[1] ? stage1[28] : stage1[26];
    assign stage2[27] = sel[1] ? stage1[29] : stage1[27];
    assign stage2[28] = sel[1] ? stage1[30] : stage1[28];
    assign stage2[29] = sel[1] ? stage1[31] : stage1[29];
    assign stage2[30] = sel[1] ? 1'b0      : stage1[30];
    assign stage2[31] = sel[1] ? 1'b0      : stage1[31];

    // Shift by 4 if sel[2] is set
    assign stage3[0]  = sel[2] ? stage2[4]  : stage2[0];
    assign stage3[1]  = sel[2] ? stage2[5]  : stage2[1];    
    assign stage3[2]  = sel[2] ? stage2[6]  : stage2[2];
    assign stage3[3]  = sel[2] ? stage2[7]  : stage2[3];
    assign stage3[4]  = sel[2] ? stage2[8]  : stage2[4];
    assign stage3[5]  = sel[2] ? stage2[9]  : stage2[5];
    assign stage3[6]  = sel[2] ? stage2[10] : stage2[6];
    assign stage3[7]  = sel[2] ? stage2[11] : stage2[7];
    assign stage3[8]  = sel[2] ? stage2[12] : stage2[8];
    assign stage3[9]  = sel[2] ? stage2[13] : stage2[9];
    assign stage3[10] = sel[2] ? stage2[14] : stage2[10];
    assign stage3[11] = sel[2] ? stage2[15] : stage2[11];
    assign stage3[12] = sel[2] ? stage2[16] : stage2[12];
    assign stage3[13] = sel[2] ? stage2[17] : stage2[13];
    assign stage3[14] = sel[2] ? stage2[18] : stage2[14];
    assign stage3[15] = sel[2] ? stage2[19] : stage2[15];
    assign stage3[16] = sel[2] ? stage2[20] : stage2[16];
    assign stage3[17] = sel[2] ? stage2[21] : stage2[17];
    assign stage3[18] = sel[2] ? stage2[22] : stage2[18];
    assign stage3[19] = sel[2] ? stage2[23] : stage2[19];
    assign stage3[20] = sel[2] ? stage2[24] : stage2[20];
    assign stage3[21] = sel[2] ? stage2[25] : stage2[21];
    assign stage3[22] = sel[2] ? stage2[26] : stage2[22];
    assign stage3[23] = sel[2] ? stage2[27] : stage2[23];
    assign stage3[24] = sel[2] ? stage2[28] : stage2[24];
    assign stage3[25] = sel[2] ? stage2[29] : stage2[25];
    assign stage3[26] = sel[2] ? stage2[30] : stage2[26];
    assign stage3[27] = sel[2] ? stage2[31] : stage2[27];
    assign stage3[28] = sel[2] ? 1'b0      : stage2[28];
    assign stage3[29] = sel[2] ? 1'b0      : stage2[29];
    assign stage3[30] = sel[2] ? 1'b0      : stage2[30];
    assign stage3[31] = sel[2] ? 1'b0      : stage2[31];
    
    // Shift by 8 if sel[3] is set
    assign stage4[0]  = sel[3] ? stage3[8]  : stage3[0];
    assign stage4[1]  = sel[3] ? stage3[9]  : stage3[1];
    assign stage4[2]  = sel[3] ? stage3[10] : stage3[2];
    assign stage4[3]  = sel[3] ? stage3[11] : stage3[3];
    assign stage4[4]  = sel[3] ? stage3[12] : stage3[4];
    assign stage4[5]  = sel[3] ? stage3[13] : stage3[5];
    assign stage4[6]  = sel[3] ? stage3[14] : stage3[6];
    assign stage4[7]  = sel[3] ? stage3[15] : stage3[7];
    assign stage4[8]  = sel[3] ? stage3[16] : stage3[8];
    assign stage4[9]  = sel[3] ? stage3[17] : stage3[9];
    assign stage4[10] = sel[3] ? stage3[18] : stage3[10];
    assign stage4[11] = sel[3] ? stage3[19] : stage3[11];
    assign stage4[12] = sel[3] ? stage3[20] : stage3[12];
    assign stage4[13] = sel[3] ? stage3[21] : stage3[13];
    assign stage4[14] = sel[3] ? stage3[22] : stage3[14];
    assign stage4[15] = sel[3] ? stage3[23] : stage3[15];
    assign stage4[16] = sel[3] ? stage3[24] : stage3[16];
    assign stage4[17] = sel[3] ? stage3[25] : stage3[17];
    assign stage4[18] = sel[3] ? stage3[26] : stage3[18];
    assign stage4[19] = sel[3] ? stage3[27] : stage3[19];
    assign stage4[20] = sel[3] ? stage3[28] : stage3[20];
    assign stage4[21] = sel[3] ? stage3[29] : stage3[21];
    assign stage4[22] = sel[3] ? stage3[30] : stage3[22];
    assign stage4[23] = sel[3] ? stage3[31] : stage3[23];
    assign stage4[24] = sel[3] ? 1'b0      : stage3[24];
    assign stage4[25] = sel[3] ? 1'b0      : stage3[25];
    assign stage4[26] = sel[3] ? 1'b0      : stage3[26];
    assign stage4[27] = sel[3] ? 1'b0      : stage3[27];
    assign stage4[28] = sel[3] ? 1'b0      : stage3[28];
    assign stage4[29] = sel[3] ? 1'b0      : stage3[29];
    assign stage4[30] = sel[3] ? 1'b0      : stage3[30];
    assign stage4[31] = sel[3] ? 1'b0      : stage3[31];

    // Shift by 16 if sel[4] is set
    assign stage5[0]  = sel[4] ? stage4[16] : stage4[0];
    assign stage5[1]  = sel[4] ? stage4[17] : stage4[1];
    assign stage5[2]  = sel[4] ? stage4[18] : stage4[2];
    assign stage5[3]  = sel[4] ? stage4[19] : stage4[3];
    assign stage5[4]  = sel[4] ? stage4[20] : stage4[4];
    assign stage5[5]  = sel[4] ? stage4[21] : stage4[5];
    assign stage5[6]  = sel[4] ? stage4[22] : stage4[6];
    assign stage5[7]  = sel[4] ? stage4[23] : stage4[7];
    assign stage5[8]  = sel[4] ? stage4[24] : stage4[8];
    assign stage5[9]  = sel[4] ? stage4[25] : stage4[9];
    assign stage5[10] = sel[4] ? stage4[26] : stage4[10];
    assign stage5[11] = sel[4] ? stage4[27] : stage4[11];
    assign stage5[12] = sel[4] ? stage4[28] : stage4[12];
    assign stage5[13] = sel[4] ? stage4[29] : stage4[13];
    assign stage5[14] = sel[4] ? stage4[30] : stage4[14];
    assign stage5[15] = sel[4] ? stage4[31] : stage4[15];
    assign stage5[16] = sel[4] ? 1'b0      : stage4[16];
    assign stage5[17] = sel[4] ? 1'b0      : stage4[17];
    assign stage5[18] = sel[4] ? 1'b0      : stage4[18];
    assign stage5[19] = sel[4] ? 1'b0      : stage4[19];
    assign stage5[20] = sel[4] ? 1'b0      : stage4[20];
    assign stage5[21] = sel[4] ? 1'b0      : stage4[21];
    assign stage5[22] = sel[4] ? 1'b0      : stage4[22];
    assign stage5[23] = sel[4] ? 1'b0      : stage4[23];
    assign stage5[24] = sel[4] ? 1'b0      : stage4[24];
    assign stage5[25] = sel[4] ? 1'b0      : stage4[25];
    assign stage5[26] = sel[4] ? 1'b0      : stage4[26];
    assign stage5[27] = sel[4] ? 1'b0      : stage4[27];
    assign stage5[28] = sel[4] ? 1'b0      : stage4[28];
    assign stage5[29] = sel[4] ? 1'b0      : stage4[29];
    assign stage5[30] = sel[4] ? 1'b0      : stage4[30];
    assign stage5[31] = sel[4] ? 1'b0      : stage4[31];

    assign y = stage2; // Final output after shifts

endmodule
